module Monster_state(clk, state);

    input wire clk;
    output reg [227: 0] state;

    always @(posedge clk) begin
        
    end

endmodule
